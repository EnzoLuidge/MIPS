library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 13;
          addrWidth: natural := 9
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is
  constant NOP  : std_logic_vector(3 downto 0) := "0000";
  constant LDA  : std_logic_vector(3 downto 0) := "0001";
  constant SOMA : std_logic_vector(3 downto 0) := "0010";
  constant SUB  : std_logic_vector(3 downto 0) := "0011";
  constant LDI : std_logic_vector(3 downto 0) := "0100";
  constant STA : std_logic_vector(3 downto 0) := "0101";
  constant JMP : std_logic_vector(3 downto 0) := "0110"; 
  constant JEQ : std_logic_vector(3 downto 0) := "0111";
  constant CEQ : std_logic_vector(3 downto 0) := "1000";
  constant JSR : std_logic_vector(3 downto 0) := "1001";
  constant RET : std_logic_vector(3 downto 0) := "1010";
  constant ANDi : std_logic_vector(3 downto 0) := "1011";
  constant ORi : std_logic_vector(3 downto 0) := "1100";
  
  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
      -- Palavra de Controle = SelMUX, Habilita_A, Reset_A, Operacao_ULA
      -- Inicializa os endereços:
tmp(0) := x"4" & '0' & x"00";	-- LDI $0  	#Carrega o acumulador com o valor 0
tmp(1) := x"5" & '1' & x"20";	-- STA @288 	#Armazena o valor do acumulador em HEX0
tmp(2) := x"5" & '1' & x"21";	-- STA @289 	#Armazena o valor do acumulador em HEX1
tmp(3) := x"5" & '1' & x"22";	-- STA @290 	#Armazena o valor do acumulador em HEX2
tmp(4) := x"5" & '1' & x"23";	-- STA @291 	#Armazena o valor do acumulador em HEX3
tmp(5) := x"5" & '1' & x"24";	-- STA @292 	#Armazena o valor do acumulador em HEX4
tmp(6) := x"5" & '1' & x"25";	-- STA @293 	#Armazena o valor do acumulador em HEX5
tmp(7) := x"0" & '0' & x"00";	-- NOP
tmp(8) := x"4" & '0' & x"00";	-- LDI $0 	#Carrega o acumulador com o valor 0
tmp(9) := x"5" & '1' & x"00";	-- STA @256 	#Armazena o valor do bit0 do acumulador no LDR0 ~ LEDR7
tmp(10) := x"5" & '1' & x"01";	-- STA @257 	#Armazena o valor do bit0 do acumulador no LDR8
tmp(11) := x"5" & '1' & x"02";	-- STA @258 	#Armazena o valor do bit0 do acumulador no LDR9
tmp(12) := x"0" & '0' & x"00";	-- NOP
tmp(13) := x"4" & '0' & x"00";	-- LDI $0 	#Carrega o acumulador com o valor 0
tmp(14) := x"5" & '0' & x"00";	-- STA @0 	#Armazena o valor do acumulador em MEM[0] unidades
tmp(15) := x"5" & '0' & x"01";	-- STA @1 	#Armazena o valor do acumulador em MEM[1] dezenas
tmp(16) := x"5" & '0' & x"02";	-- STA @2 	#Armazena o valor do acumulador em MEM[2] centenas
tmp(17) := x"5" & '0' & x"14";	-- STA @20 	#armazena o valor do acumulador em MEM[20] unidades de milhar 
tmp(18) := x"5" & '0' & x"15";	-- STA @21 	#armazena o valor do acumulador em MEM[21] dezenas de milhar
tmp(19) := x"5" & '0' & x"16";	-- STA @22 	#armazena o valor do acumulador em MEM[22] centenas de milhar
tmp(20) := x"5" & '0' & x"03";	-- STA @3 	#Armazena o valor do acumulador em MEM[3] para fazer comparacoes
tmp(21) := x"5" & '0' & x"0A";	-- STA @10 	#Armazena o valor do acumulador em MEM[10] flag de proceder com a contagem
tmp(22) := x"5" & '0' & x"3E";	-- STA @62 	#Armazena o valor do acumulador em MEM[62] flag de proceder com o decremento
tmp(23) := x"0" & '0' & x"00";	-- NOP
tmp(24) := x"4" & '0' & x"X1";	-- LDI $-1 	#Carrega o acumulador com o valor -1
tmp(25) := x"5" & '0' & x"32";	-- STA @50 	#Armazena o valor do acumulador em MEM[50] para fazer comparacao de decrementos
tmp(26) := x"4" & '0' & x"01";	-- LDI $1 	#Carrega o acumulador com o valor 1
tmp(27) := x"5" & '0' & x"04";	-- STA @4 	#Armazena o valor do acumulador em MEM[4] para fazer incrementos
tmp(28) := x"5" & '0' & x"05";	-- STA @5 	#Armazena o valor do acumulador em MEM[5] para fazer comparacoes
tmp(29) := x"5" & '1' & x"FF";	-- STA @511 	#Limpa a leitura do botão zero
tmp(30) := x"5" & '1' & x"FE";	-- STA @510 	#Limpa a leitura do botão um
tmp(31) := x"0" & '0' & x"00";	-- NOP
tmp(32) := x"4" & '0' & x"0A";	-- LDI $10 	#Carrega o acumulador com o valor 10
tmp(33) := x"5" & '0' & x"06";	-- STA @6 	#Armazena o valor do acumulador em MEM[6] para fazer comparacoes que definem o limite da faixa a ser exibida no display
tmp(34) := x"0" & '0' & x"00";	-- NOP 	#FIM DO SETUP
tmp(35) := x"9" & '0' & x"3D";	-- JSR @61
tmp(36) := x"0" & '0' & x"00";	-- NOP
tmp(37) := x"0" & '0' & x"00";	-- NOP inicio:
tmp(38) := x"1" & '1' & x"61";	-- LDA @353 	#Ler o botão de incremento de contagem KEY1 carrega o acumulador com a leitura do botão KEY1
tmp(39) := x"B" & '0' & x"05";	-- ANDi @5 	#mascara bit
tmp(40) := x"8" & '0' & x"03";	-- CEQ @3 	#Compara acumulador com o valor da memoria[3], que é 0
tmp(41) := x"7" & '0' & x"2B";	-- JEQ @43
tmp(42) := x"9" & '0' & x"92";	-- JSR @146
tmp(43) := x"0" & '0' & x"00";	-- NOP pula99:
tmp(44) := x"9" & '1' & x"12";	-- JSR @274
tmp(45) := x"0" & '0' & x"00";	-- NOP
tmp(46) := x"1" & '1' & x"60";	-- LDA @352 	#Ler/Armazenar no acumulador o botão de configuração do limite de incremento KEY1
tmp(47) := x"8" & '0' & x"03";	-- CEQ @3 	#Compara acumulador com o valor da mem[3], que é 0, ou seja, se key 1 foi pressionado
tmp(48) := x"7" & '0' & x"33";	-- JEQ @51
tmp(49) := x"9" & '0' & x"3D";	-- JSR @61
tmp(50) := x"0" & '0' & x"00";	-- NOP
tmp(51) := x"0" & '0' & x"00";	-- NOP pula98:
tmp(52) := x"9" & '0' & x"E2";	-- JSR @226
tmp(53) := x"0" & '0' & x"00";	-- NOP
tmp(54) := x"1" & '1' & x"64";	-- LDA @356 	#Ler/Armazenar o botão de reiniciar contagem FPGA_RESET
tmp(55) := x"8" & '0' & x"03";	-- CEQ @3 	# MEM[3] = 0 Caso esteja pressionado, desviar para a sub-rotina de reiniciar contagem
tmp(56) := x"7" & '0' & x"3B";	-- JEQ @59
tmp(57) := x"9" & '1' & x"06";	-- JSR @262
tmp(58) := x"0" & '0' & x"00";	-- NOP
tmp(59) := x"0" & '0' & x"00";	-- NOP pula97:
tmp(60) := x"6" & '0' & x"25";	-- JMP @37
tmp(61) := x"0" & '0' & x"00";	-- NOP limiteincremento:
tmp(62) := x"4" & '0' & x"01";	-- LDI $1
tmp(63) := x"5" & '1' & x"FF";	-- STA @511
tmp(64) := x"4" & '0' & x"01";	-- LDI $1 	#acender o led 0 indicando que iremos configurar o limite de incremento do display 0
tmp(65) := x"5" & '1' & x"00";	-- STA @256
tmp(66) := x"0" & '0' & x"00";	-- NOP loop0:
tmp(67) := x"0" & '0' & x"00";	-- NOP
tmp(68) := x"1" & '1' & x"60";	-- LDA @352 	#Aguardar o pressionamento de KEY0
tmp(69) := x"B" & '0' & x"01";	-- ANDi $1 	#mascara bit
tmp(70) := x"8" & '0' & x"03";	-- CEQ @3 	#Compara o valor do acumulador com o mem[3] que é 0
tmp(71) := x"7" & '0' & x"42";	-- JEQ @66
tmp(72) := x"0" & '0' & x"00";	-- NOP
tmp(73) := x"4" & '0' & x"01";	-- LDI $1
tmp(74) := x"5" & '1' & x"FF";	-- STA @511
tmp(75) := x"1" & '1' & x"40";	-- LDA @320 	#Ler o valor das chaves que definem o limite de contagem para as unidades
tmp(76) := x"5" & '0' & x"07";	-- STA @7 	#Armazena no mem[7] o valor do limite da contagem
tmp(77) := x"5" & '1' & x"25";	-- STA @293 	#armazena o valor das chaves em hex5 para visualizaçao do limite
tmp(78) := x"4" & '0' & x"02";	-- LDI $2 	#acender o led 1 indicando que iremos configurar o limite de incremento do display 0
tmp(79) := x"5" & '1' & x"00";	-- STA @256
tmp(80) := x"0" & '0' & x"00";	-- NOP loop1:
tmp(81) := x"0" & '0' & x"00";	-- NOP
tmp(82) := x"1" & '1' & x"60";	-- LDA @352 	#Aguardar o pressionamento de KEY0
tmp(83) := x"B" & '0' & x"01";	-- ANDi $1 	#mascara bit
tmp(84) := x"8" & '0' & x"03";	-- CEQ @3 	#compara o valor do acumulador com o mem[3] que é 0
tmp(85) := x"7" & '0' & x"50";	-- JEQ @80
tmp(86) := x"0" & '0' & x"00";	-- NOP 	#Se tiver pressionado, vai passar pelo CEQ e pelo JEQ e seguir o codigo
tmp(87) := x"5" & '1' & x"FF";	-- STA @511
tmp(88) := x"1" & '1' & x"40";	-- LDA @320 	#Ler o valor das chaves que definem o limite de contagem para as dezenas
tmp(89) := x"5" & '0' & x"08";	-- STA @8 	#Armazena no mem[8] o valor do limite da contagem
tmp(90) := x"5" & '1' & x"25";	-- STA @293 	#armazena o valor das chaves em hex5 para visualizaçao do limite
tmp(91) := x"4" & '0' & x"04";	-- LDI $4 	#acender o led 2 indicando que iremos configurar o limite de incremento do display 0
tmp(92) := x"5" & '1' & x"00";	-- STA @256
tmp(93) := x"0" & '0' & x"00";	-- NOP loop2:
tmp(94) := x"0" & '0' & x"00";	-- NOP
tmp(95) := x"1" & '1' & x"60";	-- LDA @352 	#Aguardar o pressionamento de KEY0
tmp(96) := x"B" & '0' & x"01";	-- ANDi $1 	#mascara bit
tmp(97) := x"8" & '0' & x"03";	-- CEQ @3 	#Compara o valor do acumulador com o mem[3] que é 0
tmp(98) := x"7" & '0' & x"5D";	-- JEQ @93
tmp(99) := x"0" & '0' & x"00";	-- NOP 	#se tiver pressionado, vai passar pelo ceq e pelo jeq e seguir o codigo
tmp(100) := x"5" & '1' & x"FF";	-- STA @511
tmp(101) := x"1" & '1' & x"40";	-- LDA @320 	#Ler o valor das chaves que definem o limite de contagem para as centenas
tmp(102) := x"5" & '0' & x"09";	-- STA @9 	#Armazena o valor no mem[9] o valor do limite da contagem 
tmp(103) := x"5" & '1' & x"25";	-- STA @293 	#armazena o valor das chaves em hex5 para visualizaçao do limite
tmp(104) := x"4" & '0' & x"08";	-- LDI $8 	#acender o led 3 indicando que iremos configurar o limite de incremento do display 0
tmp(105) := x"5" & '1' & x"00";	-- STA @256
tmp(106) := x"0" & '0' & x"00";	-- NOP loop3:
tmp(107) := x"0" & '0' & x"00";	-- NOP
tmp(108) := x"1" & '1' & x"60";	-- LDA @352 	#Aguardar o pressionamento de KEY0
tmp(109) := x"B" & '0' & x"01";	-- ANDi $1 	#mascara bit
tmp(110) := x"8" & '0' & x"03";	-- CEQ @3 	#Compara o valor do acumulador com o mem[3] que é 0
tmp(111) := x"7" & '0' & x"6A";	-- JEQ @106
tmp(112) := x"0" & '0' & x"00";	-- NOP 	#se tiver pressionado, vai passar pelo ceq e pelo jeq e seguir o codigo
tmp(113) := x"5" & '1' & x"FF";	-- STA @511
tmp(114) := x"1" & '1' & x"40";	-- LDA @320 	#Ler o valor das chaves que definem o limite de contagem para as unid de milhar
tmp(115) := x"5" & '0' & x"1E";	-- STA @30 	#Armazena o valor no mem[30] o valor do limite da contagem 
tmp(116) := x"5" & '1' & x"25";	-- STA @293 	#armazena o valor das chaves em hex5 para visualizaçao do limite
tmp(117) := x"4" & '0' & x"10";	-- LDI $16 	#acender o led 4 indicando que iremos configurar o limite de incremento do display 0
tmp(118) := x"5" & '1' & x"00";	-- STA @256
tmp(119) := x"0" & '0' & x"00";	-- NOP loop4:
tmp(120) := x"0" & '0' & x"00";	-- NOP
tmp(121) := x"1" & '1' & x"60";	-- LDA @352 	#Aguardar o pressionamento de KEY0
tmp(122) := x"B" & '0' & x"01";	-- ANDi $1 	#mascara bit
tmp(123) := x"8" & '0' & x"03";	-- CEQ @3 	#Compara o valor do acumulador com o mem[3] que é 0
tmp(124) := x"7" & '0' & x"77";	-- JEQ @119
tmp(125) := x"0" & '0' & x"00";	-- NOP 	#se tiver pressionado, vai passar pelo ceq e pelo jeq e seguir o codigo
tmp(126) := x"5" & '1' & x"FF";	-- STA @511
tmp(127) := x"1" & '1' & x"40";	-- LDA @320 	#Ler o valor das chaves que definem o limite de contagem para as dezenas de milhar
tmp(128) := x"5" & '0' & x"1F";	-- STA @31 	#Armazena o valor no mem[30] o valor do limite da contagem 
tmp(129) := x"5" & '1' & x"25";	-- STA @293 	#armazena o valor das chaves em hex5 para visualizaçao do limite
tmp(130) := x"4" & '0' & x"20";	-- LDI $32 	#acender o led 5 indicando que iremos configurar o limite de incremento do display 0
tmp(131) := x"5" & '1' & x"00";	-- STA @256
tmp(132) := x"0" & '0' & x"00";	-- NOP loop5:
tmp(133) := x"0" & '0' & x"00";	-- NOP
tmp(134) := x"1" & '1' & x"60";	-- LDA @352 	#Aguardar o pressionamento de KEY0
tmp(135) := x"B" & '0' & x"01";	-- ANDi $1 	#mascara bit
tmp(136) := x"8" & '0' & x"03";	-- CEQ @3 	#Compara o valor do acumulador com o mem[3] que é 0
tmp(137) := x"7" & '0' & x"84";	-- JEQ @132
tmp(138) := x"0" & '0' & x"00";	-- NOP 	#se tiver pressionado, vai passar pelo ceq e pelo jeq e seguir o codigo
tmp(139) := x"5" & '1' & x"FF";	-- STA @511
tmp(140) := x"1" & '1' & x"40";	-- LDA @320 	#Ler o valor das chaves que definem o limite de contagem para as centenas de milhar
tmp(141) := x"5" & '0' & x"20";	-- STA @32 	#Armazena o valor no mem[32] o valor do limite da contagem 
tmp(142) := x"5" & '1' & x"25";	-- STA @293 	#armazena o valor das chaves em hex5 para visualizaçao do limite
tmp(143) := x"4" & '0' & x"00";	-- LDI $0 	#apagar o led 
tmp(144) := x"5" & '1' & x"00";	-- STA @256
tmp(145) := x"A" & '0' & x"00";	-- RET 	#Retornar para o inicio
tmp(146) := x"0" & '0' & x"00";	-- NOP incremento:
tmp(147) := x"5" & '1' & x"FE";	-- STA @510 	#Limpar o _flag_ de botão 0 apertado acessar endereço 511.
tmp(148) := x"4" & '0' & x"00";	-- LDI $0 	#Verificar _FLAG_ de proceder com a contagem
tmp(149) := x"8" & '0' & x"0A";	-- CEQ @10 	#se estiver setado, retornar da sub rotina
tmp(150) := x"7" & '0' & x"98";	-- JEQ @152
tmp(151) := x"A" & '0' & x"00";	-- RET 	#retorno da sub rotina de jeq
tmp(152) := x"0" & '0' & x"00";	-- NOP incrementaunidade:
tmp(153) := x"4" & '0' & x"01";	-- LDI $1 	#incrementar o valor de unidades da contagem
tmp(154) := x"2" & '0' & x"00";	-- SOMA @0 	#incremento do acumulador com 1 e da mem[0], que é o valor das unidades 
tmp(155) := x"5" & '0' & x"0B";	-- STA @11 	#guardar o resultado da soma em mem[11], para ser usado posteriormente
tmp(156) := x"8" & '0' & x"06";	-- CEQ @6 	#compara o resultado do incremento das unidades com dez, que esta em mem[6] 
tmp(157) := x"7" & '0' & x"A1";	-- JEQ @161
tmp(158) := x"1" & '0' & x"0B";	-- LDA @11 	#se nao for igual, escreve o valor incrementado nas unidades
tmp(159) := x"5" & '0' & x"00";	-- STA @0 	#armazena no valor das unidades 
tmp(160) := x"A" & '0' & x"00";	-- RET 	#retorno da sub rotina jeq
tmp(161) := x"0" & '0' & x"00";	-- NOP incrementadezena:
tmp(162) := x"4" & '0' & x"00";	-- LDI $0 	#se for igual..
tmp(163) := x"5" & '0' & x"00";	-- STA @0 	#armazena 0 nas unidades 
tmp(164) := x"4" & '0' & x"01";	-- LDI $1
tmp(165) := x"2" & '0' & x"01";	-- SOMA @1 	#soma 1 do acumulador com mem[1], que é das dezenas
tmp(166) := x"5" & '0' & x"0B";	-- STA @11 	#guarda o resultado da soma em mem[11], para ser usado posteriormente 
tmp(167) := x"8" & '0' & x"06";	-- CEQ @6 	#comparando as dezenas com mem[6], que é 10
tmp(168) := x"7" & '0' & x"AD";	-- JEQ @173
tmp(169) := x"0" & '0' & x"00";	-- NOP 	#se não for igual, armazena o resultado em mem[1] das dezenas
tmp(170) := x"1" & '0' & x"0B";	-- LDA @11 
tmp(171) := x"5" & '0' & x"01";	-- STA @1 	#armazena o resultado em mem[1], das dezenas 
tmp(172) := x"A" & '0' & x"00";	-- RET 	#retorno da sub rotina jeq
tmp(173) := x"0" & '0' & x"00";	-- NOP incrementacentena:
tmp(174) := x"4" & '0' & x"00";	-- LDI $0 	#se for igual..
tmp(175) := x"5" & '0' & x"01";	-- STA @1 	#escreve 0 nas dezenas  
tmp(176) := x"4" & '0' & x"01";	-- LDI $1
tmp(177) := x"2" & '0' & x"02";	-- SOMA @2 	#soma 1 do acumulador com mem[2] que é das centenas 
tmp(178) := x"5" & '0' & x"0B";	-- STA @11 	#guarda o resultado da soma em mem[11], para ser usado posteriormente
tmp(179) := x"8" & '0' & x"06";	-- CEQ @6 	#compara as centenas com mem[6], que é 10
tmp(180) := x"7" & '0' & x"B9";	-- JEQ @185
tmp(181) := x"0" & '0' & x"00";	-- NOP 	#fim das comparações das dezenas com 10
tmp(182) := x"1" & '0' & x"0B";	-- LDA @11
tmp(183) := x"5" & '0' & x"02";	-- STA @2 	#armazena em centenas 
tmp(184) := x"A" & '0' & x"00";	-- RET 	#retorno da sub rotina jeq
tmp(185) := x"0" & '0' & x"00";	-- NOP incrementaunidadedemilhar:
tmp(186) := x"4" & '0' & x"00";	-- LDI $0 	#se for igual..
tmp(187) := x"5" & '0' & x"02";	-- STA @2 	#armazena 0 nas centenas 
tmp(188) := x"4" & '0' & x"01";	-- LDI $1
tmp(189) := x"2" & '0' & x"14";	-- SOMA @20 	#soma 1 do acumulador com mem[20], que é das unid de milhar
tmp(190) := x"5" & '0' & x"0B";	-- STA @11 	#guarda o resultado da soma em mem[11], para ser usado posteriormente 
tmp(191) := x"8" & '0' & x"06";	-- CEQ @6 	#comparando as dezenas com mem[6], que é 10
tmp(192) := x"7" & '0' & x"C5";	-- JEQ @197
tmp(193) := x"0" & '0' & x"00";	-- NOP 	#se não for igual, armazena o resultado em mem[1] das dezenas
tmp(194) := x"1" & '0' & x"0B";	-- LDA @11 
tmp(195) := x"5" & '0' & x"14";	-- STA @20 	#armazena o resultado em mem[20], das unidades de milhar 
tmp(196) := x"A" & '0' & x"00";	-- RET 	#retorno da sub rotina jeq
tmp(197) := x"0" & '0' & x"00";	-- NOP incrementadezenademilhar:
tmp(198) := x"4" & '0' & x"00";	-- LDI $0 	#se for igual..
tmp(199) := x"5" & '0' & x"14";	-- STA @20 	#armazena 0 nas unidades de milhar 
tmp(200) := x"4" & '0' & x"01";	-- LDI $1
tmp(201) := x"2" & '0' & x"15";	-- SOMA @21 	#soma 1 do acumulador com mem[21], que é das dezenas de milhar
tmp(202) := x"5" & '0' & x"0B";	-- STA @11 	#guarda o resultado da soma em mem[11], para ser usado posteriormente 
tmp(203) := x"8" & '0' & x"06";	-- CEQ @6 	#comparando as dezenas com mem[6], que é 10
tmp(204) := x"7" & '0' & x"D1";	-- JEQ @209
tmp(205) := x"0" & '0' & x"00";	-- NOP 	#se não for igual, armazena o resultado em mem[1] das dezenas
tmp(206) := x"1" & '0' & x"0B";	-- LDA @11 
tmp(207) := x"5" & '0' & x"15";	-- STA @21 	#armazena o resultado em mem[20], das dezenas de milhar 
tmp(208) := x"A" & '0' & x"00";	-- RET 	#retorno da sub rotina jeq
tmp(209) := x"0" & '0' & x"00";	-- NOP incrementacentenademilhar:
tmp(210) := x"4" & '0' & x"00";	-- LDI $0 	#se for igual..
tmp(211) := x"5" & '0' & x"15";	-- STA @21 	#armazena 0 nas unidades de milhar 
tmp(212) := x"4" & '0' & x"01";	-- LDI $1
tmp(213) := x"2" & '0' & x"16";	-- SOMA @22 	#soma 1 do acumulador com mem[22], que é das centenas de milhar
tmp(214) := x"5" & '0' & x"0B";	-- STA @11 	#guarda o resultado da soma em mem[11], para ser usado posteriormente 
tmp(215) := x"8" & '0' & x"06";	-- CEQ @6 	#comparando as dezenas com mem[6], que é 10
tmp(216) := x"7" & '0' & x"DD";	-- JEQ @221
tmp(217) := x"0" & '0' & x"00";	-- NOP 	#se não for igual, armazena o resultado em mem[1] das dezenas
tmp(218) := x"1" & '0' & x"0B";	-- LDA @11 
tmp(219) := x"5" & '0' & x"16";	-- STA @22 	#armazena o resultado em mem[22], das centenas de milhar 
tmp(220) := x"A" & '0' & x"00";	-- RET 	#retorno da sub rotina jeq
tmp(221) := x"0" & '0' & x"00";	-- NOP pula3:
tmp(222) := x"4" & '0' & x"01";	-- LDI $1 
tmp(223) := x"5" & '1' & x"01";	-- STA @257 	#led indicador de overflow LED8
tmp(224) := x"5" & '0' & x"0A";	-- STA @10 	#ativar flag de inibir contagem
tmp(225) := x"A" & '0' & x"00";	-- RET 	#retorno da sub rotina jeq
tmp(226) := x"0" & '0' & x"00";	-- NOP limitecontagem:
tmp(227) := x"1" & '0' & x"07";	-- LDA @7  	#para as unidades 
tmp(228) := x"8" & '0' & x"00";	-- CEQ @0 	#compara limite de contagem mem[7], que é das unidades, com mem[0], que é unidades 
tmp(229) := x"7" & '0' & x"E7";	-- JEQ @231
tmp(230) := x"A" & '0' & x"00";	-- RET 	#se nao for igual, retorna
tmp(231) := x"0" & '0' & x"00";	-- NOP pula4:
tmp(232) := x"1" & '0' & x"08";	-- LDA @8 	#para as dezenas 
tmp(233) := x"8" & '0' & x"01";	-- CEQ @1 	#compara limite de contagem mem[8], que é das dezenas, com mem[1], que é dezenas 
tmp(234) := x"7" & '0' & x"EC";	-- JEQ @236
tmp(235) := x"A" & '0' & x"00";	-- RET 	#se nao for igual, retorna
tmp(236) := x"0" & '0' & x"00";	-- NOP pula5:
tmp(237) := x"1" & '0' & x"09";	-- LDA @9 	#para as centenas 
tmp(238) := x"8" & '0' & x"02";	-- CEQ @2 	#compara limite de contagem mem[9], que é das centenas, com mem[2], que é centenas
tmp(239) := x"7" & '0' & x"F1";	-- JEQ @241
tmp(240) := x"A" & '0' & x"00";	-- RET 	#se nao for igual, retorna
tmp(241) := x"0" & '0' & x"00";	-- NOP pula6:
tmp(242) := x"1" & '0' & x"1E";	-- LDA @30 	#para as unid de milhar 
tmp(243) := x"8" & '0' & x"14";	-- CEQ @20 	#compara limite de contagem mem[9], que é das centenas, com mem[2], que é unid de milhar
tmp(244) := x"7" & '0' & x"F6";	-- JEQ @246
tmp(245) := x"A" & '0' & x"00";	-- RET 	#se nao for igual, retorna
tmp(246) := x"0" & '0' & x"00";	-- NOP pula7:
tmp(247) := x"1" & '0' & x"1F";	-- LDA @31 	#para as dezenas de milhar 
tmp(248) := x"8" & '0' & x"15";	-- CEQ @21 	#compara limite de contagem mem[9], que é das centenas, com mem[2], que é centenas
tmp(249) := x"7" & '0' & x"FB";	-- JEQ @251
tmp(250) := x"A" & '0' & x"00";	-- RET 	#se nao for igual, retorna
tmp(251) := x"0" & '0' & x"00";	-- NOP pula8:
tmp(252) := x"1" & '0' & x"20";	-- LDA @32 	#para as centenas de milhar
tmp(253) := x"8" & '0' & x"16";	-- CEQ @22 	#compara limite de contagem mem[9], que é das centenas, com mem[2], que é centenas
tmp(254) := x"7" & '1' & x"00";	-- JEQ @256
tmp(255) := x"A" & '0' & x"00";	-- RET 	#se nao for igual, retorna
tmp(256) := x"0" & '0' & x"00";	-- NOP pula9:
tmp(257) := x"4" & '0' & x"01";	-- LDI $1 	#ativa a flag de inibir contagem
tmp(258) := x"5" & '0' & x"0A";	-- STA @10 
tmp(259) := x"5" & '1' & x"02";	-- STA @258 	#acende o led de limite atingido LED9
tmp(260) := x"0" & '0' & x"00";	-- NOP 
tmp(261) := x"A" & '0' & x"00";	-- RET    	#retorno da sub rotina jeq
tmp(262) := x"0" & '0' & x"00";	-- NOP reinicio:
tmp(263) := x"4" & '0' & x"00";	-- LDI $0 	#escrever zero nas variaveis de contagem 
tmp(264) := x"5" & '0' & x"00";	-- STA @0 
tmp(265) := x"5" & '0' & x"01";	-- STA @1 
tmp(266) := x"5" & '0' & x"02";	-- STA @2 
tmp(267) := x"5" & '0' & x"0A";	-- STA @10 	#limpar o flag de inibir contagem
tmp(268) := x"5" & '1' & x"01";	-- STA @257 	#apagar led de overflow
tmp(269) := x"5" & '1' & x"02";	-- STA @258 	#apagar led de limite atingido
tmp(270) := x"4" & '0' & x"01";	-- LDI $1
tmp(271) := x"5" & '1' & x"FF";	-- STA @511 	#limpar key0
tmp(272) := x"5" & '1' & x"FE";	-- STA @510 	#limpar key1
tmp(273) := x"A" & '0' & x"00";	-- RET 	#retorno da sub rotina
tmp(274) := x"0" & '0' & x"00";	-- NOP escrevedisplay:
tmp(275) := x"1" & '0' & x"00";	-- LDA @0 	#armazena o valor de mem[0], das unidades, no display 
tmp(276) := x"5" & '1' & x"20";	-- STA @288
tmp(277) := x"1" & '0' & x"01";	-- LDA @1 	#armazena o valor de mem[1], das dezenas, no display 
tmp(278) := x"5" & '1' & x"21";	-- STA @289 
tmp(279) := x"1" & '0' & x"02";	-- LDA @2 	#armazena o valor de mem[2], das centenas, no display 
tmp(280) := x"5" & '1' & x"22";	-- STA @290
tmp(281) := x"1" & '0' & x"14";	-- LDA @20 	#armazena o valor de mem[20], das unidades de milhar, no display 
tmp(282) := x"5" & '1' & x"23";	-- STA @291
tmp(283) := x"1" & '0' & x"15";	-- LDA @21 	#armazena o valor de mem[21], das dezenas de milhar, no display 
tmp(284) := x"5" & '1' & x"24";	-- STA @292
tmp(285) := x"1" & '0' & x"16";	-- LDA @22 	#armazena o valor de mem[22], das centenas de milhar, no display 
tmp(286) := x"5" & '1' & x"25";	-- STA @293
tmp(287) := x"0" & '0' & x"00";	-- NOP decremento:
tmp(288) := x"5" & '1' & x"FD";	-- STA @509 	# Limpar o _flag_ de botão 0 apertado acessar endereço 511
tmp(289) := x"1" & '0' & x"00";	-- LDA @0     	# Carregar valor das unidades
tmp(290) := x"8" & '0' & x"00";	-- CEQ @0     	# Verificar se as unidades são zero
tmp(291) := x"7" & '1' & x"26";	-- JEQ @294
tmp(292) := x"4" & '0' & x"01";	-- LDI $1     	# Se as unidades não forem zero, continuar com o decremento
tmp(293) := x"6" & '1' & x"45";	-- JMP @325
tmp(294) := x"0" & '0' & x"00";	-- NOP verificaDezena:
tmp(295) := x"1" & '0' & x"01";	-- LDA @1     	# Carregar valor das dezenas
tmp(296) := x"8" & '0' & x"00";	-- CEQ @0     	# Verificar se as dezenas são zero
tmp(297) := x"7" & '1' & x"2C";	-- JEQ @300
tmp(298) := x"4" & '0' & x"01";	-- LDI $1     	# Se as dezenas não forem zero, continuar com o decremento
tmp(299) := x"6" & '1' & x"45";	-- JMP @325
tmp(300) := x"0" & '0' & x"00";	-- NOP verificaCentena:
tmp(301) := x"1" & '0' & x"02";	-- LDA @2     	# Carregar valor das centenas
tmp(302) := x"8" & '0' & x"00";	-- CEQ @0     	# Verificar se as centenas são zero
tmp(303) := x"7" & '1' & x"32";	-- JEQ @306
tmp(304) := x"4" & '0' & x"01";	-- LDI $1     	# Se as centenas não forem zero, continuar com o decremento
tmp(305) := x"6" & '1' & x"45";	-- JMP @325
tmp(306) := x"0" & '0' & x"00";	-- NOP verificaUnidadeMilhar:
tmp(307) := x"1" & '0' & x"14";	-- LDA @20    	# Carregar valor das unidades de milhar
tmp(308) := x"8" & '0' & x"00";	-- CEQ @0     	# Verificar se as unidades de milhar são zero
tmp(309) := x"7" & '1' & x"38";	-- JEQ @312
tmp(310) := x"4" & '0' & x"01";	-- LDI $1     	# Se as unidades de milhar não forem zero, continuar com o decremento
tmp(311) := x"6" & '1' & x"45";	-- JMP @325
tmp(312) := x"0" & '0' & x"00";	-- NOP verificaDezenaMilhar:
tmp(313) := x"1" & '0' & x"15";	-- LDA @21    	# Carregar valor das dezenas de milhar
tmp(314) := x"8" & '0' & x"00";	-- CEQ @0     	# Verificar se as dezenas de milhar são zero
tmp(315) := x"7" & '1' & x"3E";	-- JEQ @318
tmp(316) := x"4" & '0' & x"01";	-- LDI $1     	# Se as dezenas de milhar não forem zero, continuar com o decremento
tmp(317) := x"6" & '1' & x"45";	-- JMP @325
tmp(318) := x"0" & '0' & x"00";	-- NOP verificaCentenaMilhar:
tmp(319) := x"1" & '0' & x"16";	-- LDA @22    	# Carregar valor das centenas de milhar
tmp(320) := x"8" & '0' & x"00";	-- CEQ @0     	# Verificar se as centenas de milhar são zero
tmp(321) := x"7" & '1' & x"81";	-- JEQ @385
tmp(322) := x"4" & '0' & x"01";	-- LDI $1     	# Se as centenas de milhar não forem zero, continuar com o decremento
tmp(323) := x"7" & '1' & x"45";	-- JEQ @325
tmp(324) := x"A" & '0' & x"00";	-- RET 	# Retorno da sub-rotina de jeq
tmp(325) := x"0" & '0' & x"00";	-- NOP decrementacentenademilhar:
tmp(326) := x"4" & '0' & x"01";	-- LDI $1 	# Decrementar o valor das centenas de milhar da contagem
tmp(327) := x"3" & '0' & x"16";	-- SUB @22 	# Subtrair 1 do acumulador com mem[22], que é das centenas de milhar
tmp(328) := x"5" & '0' & x"0B";	-- STA @11 	# Guardar o resultado da subtração em mem[11], para ser usado posteriormente
tmp(329) := x"8" & '0' & x"32";	-- CEQ @50 	# Comparar o resultado da subtração das centenas de milhar com -1
tmp(330) := x"7" & '1' & x"4F";	-- JEQ @335
tmp(331) := x"0" & '0' & x"00";	-- NOP 	# Se não for igual, armazenar o resultado em mem[22] das centenas de milhar
tmp(332) := x"1" & '0' & x"0B";	-- LDA @11 
tmp(333) := x"5" & '0' & x"16";	-- STA @22 	# Armazenar o resultado em mem[22], das centenas de milhar
tmp(334) := x"A" & '0' & x"00";	-- RET 	# Retorno da sub-rotina de jeq
tmp(335) := x"0" & '0' & x"00";	-- NOP decrementadezenademilhar:
tmp(336) := x"4" & '0' & x"01";	-- LDI $1 	# Decrementar o valor das dezenas de milhar da contagem
tmp(337) := x"3" & '0' & x"15";	-- SUB @21 	# Subtrair 1 do acumulador com mem[21], que é das dezenas de milhar
tmp(338) := x"5" & '0' & x"0B";	-- STA @11 	# Guardar o resultado da subtração em mem[11], para ser usado posteriormente
tmp(339) := x"8" & '0' & x"32";	-- CEQ @50 	# Comparar o resultado da subtração das dezenas de milhar com -1
tmp(340) := x"7" & '1' & x"59";	-- JEQ @345
tmp(341) := x"0" & '0' & x"00";	-- NOP 	# Se não for igual, armazenar o resultado em mem[21] das dezenas de milhar
tmp(342) := x"1" & '0' & x"0B";	-- LDA @11 
tmp(343) := x"5" & '0' & x"15";	-- STA @21 	# Armazenar o resultado em mem[21], das dezenas de milhar
tmp(344) := x"A" & '0' & x"00";	-- RET 	# Retorno da sub-rotina de jeq
tmp(345) := x"0" & '0' & x"00";	-- NOP decrementaunidadedemilhar:
tmp(346) := x"4" & '0' & x"01";	-- LDI $1 	# Decrementar o valor das unidades de milhar da contagem
tmp(347) := x"3" & '0' & x"14";	-- SUB @20 	# Subtrair 1 do acumulador com mem[20], que é das unidades de milhar
tmp(348) := x"5" & '0' & x"0B";	-- STA @11 	# Guardar o resultado da subtração em mem[11], para ser usado posteriormente
tmp(349) := x"8" & '0' & x"32";	-- CEQ @50 	# Comparar o resultado da subtração das unidades de milhar com -1
tmp(350) := x"7" & '1' & x"63";	-- JEQ @355
tmp(351) := x"0" & '0' & x"00";	-- NOP 	# Se não for igual, armazenar o resultado em mem[20] das unidades de milhar
tmp(352) := x"1" & '0' & x"0B";	-- LDA @11 
tmp(353) := x"5" & '0' & x"14";	-- STA @20 	# Armazenar o resultado em mem[20], das unidades de milhar
tmp(354) := x"A" & '0' & x"00";	-- RET 	# Retorno da sub-rotina de jeq
tmp(355) := x"0" & '0' & x"00";	-- NOP decrementacentena:
tmp(356) := x"4" & '0' & x"01";	-- LDI $1 	# Decrementar o valor das centenas da contagem
tmp(357) := x"3" & '0' & x"02";	-- SUB @2 	# Subtrair 1 do acumulador com mem[2], que é das centenas
tmp(358) := x"5" & '0' & x"0B";	-- STA @11 	# Guardar o resultado da subtração em mem[11], para ser usado posteriormente
tmp(359) := x"8" & '0' & x"32";	-- CEQ @50 	# Comparar o resultado da subtração das centenas com -1
tmp(360) := x"7" & '1' & x"6D";	-- JEQ @365
tmp(361) := x"0" & '0' & x"00";	-- NOP 	# Se não for igual, armazenar o resultado em mem[2] das centenas
tmp(362) := x"1" & '0' & x"0B";	-- LDA @11 
tmp(363) := x"5" & '0' & x"02";	-- STA @2 	# Armazenar o resultado em mem[2], das centenas
tmp(364) := x"A" & '0' & x"00";	-- RET 	# Retorno da sub-rotina de jeq
tmp(365) := x"0" & '0' & x"00";	-- NOP decrementadezena:
tmp(366) := x"4" & '0' & x"01";	-- LDI $1 	# Decrementar o valor das dezenas da contagem
tmp(367) := x"3" & '0' & x"01";	-- SUB @1 	# Subtrair 1 do acumulador com mem[1], que é das dezenas
tmp(368) := x"5" & '0' & x"0B";	-- STA @11 	# Guardar o resultado da subtração em mem[11], para ser usado posteriormente
tmp(369) := x"8" & '0' & x"32";	-- CEQ @50 	# Comparar o resultado da subtração das dezenas com -1
tmp(370) := x"7" & '1' & x"77";	-- JEQ @375
tmp(371) := x"0" & '0' & x"00";	-- NOP 	# Se não for igual, armazenar o resultado em mem[1] das dezenas
tmp(372) := x"1" & '0' & x"0B";	-- LDA @11 
tmp(373) := x"5" & '0' & x"01";	-- STA @1 	# Armazenar o resultado em mem[1], das dezenas
tmp(374) := x"A" & '0' & x"00";	-- RET 	# Retorno da sub-rotina de jeq
tmp(375) := x"0" & '0' & x"00";	-- NOP decrementaunidade:
tmp(376) := x"4" & '0' & x"01";	-- LDI $1 	# Decrementar o valor das unidades da contagem
tmp(377) := x"3" & '0' & x"00";	-- SUB @0 	# Subtrair 1 do acumulador com mem[0], que é das unidades
tmp(378) := x"5" & '0' & x"0B";	-- STA @11 	# Guardar o resultado da subtração em mem[11], para ser usado posteriormente
tmp(379) := x"8" & '0' & x"32";	-- CEQ @50 	# Comparar o resultado da subtração das unidades com -1
tmp(380) := x"7" & '1' & x"81";	-- JEQ @385
tmp(381) := x"0" & '0' & x"00";	-- NOP 	# Se não for igual, armazenar o resultado em mem[0] das unidades
tmp(382) := x"1" & '0' & x"0B";	-- LDA @11 
tmp(383) := x"5" & '0' & x"00";	-- STA @0 	# Armazenar o resultado em mem[0], das unidades
tmp(384) := x"A" & '0' & x"00";	-- RET 	# Retorno da sub-rotina de jeq
tmp(385) := x"0" & '0' & x"00";	-- NOP pula15:
tmp(386) := x"4" & '0' & x"02";	-- LDI $2
tmp(387) := x"5" & '1' & x"02";	-- STA @258 	# led indicador de limite atingido LED8
tmp(388) := x"A" & '0' & x"00";	-- RET 	# Retorno da sub-rotina jeq

        return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;